module OR(A, B, F);
    input[7:0] A, B;
    output[7:0] F;
    assign F = A | B;
endmodule